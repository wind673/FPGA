`timescale 1ns/1ps
module LED_Test;
reg clk; 
reg rst_n;
wire [3:0] led ;

initial 
	begin
		clk = 1;
		rst_n = 0;
		#20.1
		rst_n = 1;
		#20000
		$stop ;
	end
always #10 clk <= ~clk ;
LED Test1 (
    .clk(clk), // 开发板上输入时钟: 50Mhz
    .rst_n(rst_n), // 开发板上输入复位按键
    .led (led)// 输出 LED 灯,用于控制开发板上四个 LED(LED1~LED4)
);



endmodule 



