library verilog;
use verilog.vl_types.all;
entity LED_vlg_tst is
end LED_vlg_tst;
